module core(
	input wire clk,
	input wire [31:0]  datain0, datain1, datain2, datain3,
	output wire [31:0] dataout0, dataout1, dataout2, dataout3
);
	
	endmodule